* Extracted by KLayout with SG13G2 LVS runset on : 01/09/2025 07:07

.SUBCKT M34 PQ XY YX
M$1 XY YX PQ \$3 sg13_lv_nmos L=0.13u W=8u AS=2.12p AD=2.12p PS=16.24u PD=16.24u
.ENDS M34
