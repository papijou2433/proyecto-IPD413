** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/proyecto-IPD413/klayout/LVS/M7.sch
.subckt M7

M1 Vss CLK common Vss sg13_lv_nmos l=0.13u w=1.0u ng=1 m=15
.ends
.end
