** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/proyecto-IPD413/klayout/LVS/M12.sch
.subckt M12

M1 common Vin12 PQ Vss sg13_lv_nmos l=0.5u w=2.5u ng=5 m=8
.ends
.end
