* Extracted by KLayout with SG13G2 LVS runset on : 01/09/2025 03:52

.SUBCKT M89 Vdd CLK PQ
M$1 Vdd CLK PQ Vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=5.36u PD=5.36u
.ENDS M89
