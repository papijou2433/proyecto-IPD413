* Extracted by KLayout with SG13G2 LVS runset on : 01/09/2025 02:24

.SUBCKT M7
X$1 \$1 \$4 \$2 \$3 \$I3 M7_row
X$2 \$1 \$4 \$2 \$3 \$I3 M7_row
X$3 \$1 \$4 \$2 \$3 \$I3 M7_row
.ENDS M7

.SUBCKT M7_row \$1 \$I12 \$I11 \$I9 \$I8
X$1 \$1 \$I8 \$I12 M7_single
X$2 \$1 \$I8 \$I11 M7_single
X$3 \$1 \$I8 \$I11 M7_single
X$4 \$1 \$I8 \$I9 M7_single
X$5 \$1 \$I8 \$I9 M7_single
.ENDS M7_row

.SUBCKT M7_single \$1 \$2 \$3
X$1 \$1 \$3 \$1 \$2 nmos
.ENDS M7_single

.SUBCKT nmos \$1 \$2 \$3 \$5
M$1 \$1 \$5 \$2 \$3 sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
.ENDS nmos
