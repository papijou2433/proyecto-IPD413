** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/proyecto-IPD413/xschem/TB/TB_lvPMOS_cgate-ext.sch
.subckt TB_lvPMOS_cgate-ext

R1 VOUT VIN 1k m=1
V1 VIN GND PULSE (1 0 0 1p 1p {T/2} {T})
V1V V1V GND 1
R2 VOUT_C VIN_C 1k m=1
V2 VIN_C GND PULSE (1 0 0 1p 1p {T/2} {T})
C1 V1V VOUT_C {Co} m=1
M1 V1V VOUT V1V V1V sg13_lv_pmos w=1.0u l=0.13u ng=1 m=1
**** begin user architecture code



.param T = 1.6u
.param Co = 119.8p
.tran 10p {T}
.save all
.ic v(vout) = 1
.control
run
meas tran teval WHEN v(vout) = 0.37
let res_val = 1000
let cap_val = teval/res_val
plot v(vin) v(vout) v(vout_c)
print cap_val
.endc




.lib cornerMOShv.lib mos_tt
.lib cornerMOSlv.lib mos_tt
*.lib cornerMOShv.lib mos_ff
*.lib cornerMOSlv.lib mos_ff
*.lib cornerMOShv.lib mos_ss
*.lib cornerMOSlv.lib mos_ss
*.lib cornerMOShv.lib mos_sf
*.lib cornerMOSlv.lib mos_sf
*.lib cornerMOShv.lib mos_fs
*.lib cornerMOSlv.lib mos_fs

.include /opt/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ
*.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/diodes.lib



*M1 hvPMOS
.param temp=27
.param mult_M1 = 12000
.param w_M1 =10u
.param l_M1 = 0.4u
.param ng_M1 = 1

*M2 hvNMOS
.param mult_M2 = 4000
.param w_M2 =10u
.param l_M2 =0.45u
.param ng_M2 =1






**** end user architecture code
.ends
.GLOBAL GND
.end
